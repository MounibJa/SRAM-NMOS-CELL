magic
tech sky130A
magscale 1 2
timestamp 1764459837
<< nmos >>
rect -25 -45 25 45
<< ndiff >>
rect -83 33 -25 45
rect -83 -33 -71 33
rect -37 -33 -25 33
rect -83 -45 -25 -33
rect 25 33 83 45
rect 25 -33 37 33
rect 71 -33 83 33
rect 25 -45 83 -33
<< ndiffc >>
rect -71 -33 -37 33
rect 37 -33 71 33
<< poly >>
rect -33 117 33 133
rect -33 83 -17 117
rect 17 83 33 117
rect -33 67 33 83
rect -25 45 25 67
rect -25 -67 25 -45
rect -33 -83 33 -67
rect -33 -117 -17 -83
rect 17 -117 33 -83
rect -33 -133 33 -117
<< polycont >>
rect -17 83 17 117
rect -17 -117 17 -83
<< locali >>
rect -54 83 -17 117
rect 17 83 54 117
rect -71 33 -37 49
rect -71 -49 -37 -33
rect 37 33 71 49
rect 37 -49 71 -33
rect -54 -117 -17 -83
rect 17 -117 54 -83
<< viali >>
rect -17 83 17 117
rect -71 -33 -37 33
rect 37 -33 71 33
rect -17 -117 17 -83
<< metal1 >>
rect -29 117 29 123
rect -54 83 -17 117
rect 17 83 54 117
rect -29 77 29 83
rect -77 33 -31 45
rect -77 -33 -71 33
rect -37 -33 -31 33
rect -77 -45 -31 -33
rect 31 33 77 45
rect 31 -33 37 33
rect 71 -33 77 33
rect 31 -45 77 -33
rect -63 -83 57 -73
rect -63 -93 -17 -83
rect 17 -93 57 -83
rect -63 -153 -23 -93
rect 37 -153 57 -93
rect -63 -173 57 -153
<< via1 >>
rect -23 -117 -17 -93
rect -17 -117 17 -93
rect 17 -117 37 -93
rect -23 -153 37 -117
<< metal2 >>
rect -43 -93 57 -73
rect -43 -153 -23 -93
rect 37 -153 57 -93
rect -43 -173 57 -153
<< labels >>
rlabel ndiffc -54 0 -54 0 0 D
port 1 nsew
rlabel ndiffc 54 0 54 0 0 S
port 2 nsew
rlabel polycont 0 100 0 100 0 G
port 3 nsew
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.450 l 0.250 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
