* NGSPICE file created from BitCellNoResis.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_BHJCXL D0 G0 S1 G1 a_79_n50# VSUBS
X0 a_79_n50# G1 S1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.25
X1 S1 G0 D0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.25
C0 a_79_n50# G1 0.00663f
C1 S1 G1 0.00663f
C2 S1 D0 0.06743f
C3 S1 G0 0.00663f
C4 a_79_n50# S1 0.06743f
C5 G1 G0 0.0147f
C6 D0 G0 0.00663f
C7 S1 VSUBS 0.03655f
C8 D0 VSUBS 0.07653f
C9 G0 VSUBS 0.21316f
C10 G1 VSUBS 0.21316f
C11 a_79_n50# VSUBS 0.07653f
.ends

.subckt sky130_fd_pr__nfet_01v8_HKHAX8 D S G VSUBS
X0 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.25
C0 G D 0.04837f
C1 G S 0.04837f
C2 D S 0.09984f
C3 S VSUBS 0.0829f
C4 D VSUBS 0.0829f
C5 G VSUBS 0.35917f
.ends

.subckt sky130_fd_pr__pfet_01v8_6KFL8S B D S G VSUBS
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=1.2
C0 B G 0.56403f
C1 B S 0.04171f
C2 B D 0.04171f
C3 S G 0.05151f
C4 G D 0.05151f
C5 S D 0.02073f
C6 S VSUBS 0.02575f
C7 D VSUBS 0.02575f
C8 G VSUBS 0.3744f
C9 B VSUBS 1.40766f
.ends

.subckt BitCellNoResis VDD GND WL BL BL_N BL_IN BL_NIN
Xsky130_fd_pr__nfet_01v8_BHJCXL_0 BL_IN BL_NIN GND BL_IN BL_NIN GND sky130_fd_pr__nfet_01v8_BHJCXL
Xsky130_fd_pr__nfet_01v8_HKHAX8_0 BL_N BL_NIN WL GND sky130_fd_pr__nfet_01v8_HKHAX8
Xsky130_fd_pr__nfet_01v8_HKHAX8_1 BL_IN BL WL GND sky130_fd_pr__nfet_01v8_HKHAX8
Xsky130_fd_pr__pfet_01v8_6KFL8S_0 VDD VDD BL_IN GND GND sky130_fd_pr__pfet_01v8_6KFL8S
Xsky130_fd_pr__pfet_01v8_6KFL8S_1 VDD BL_NIN VDD GND GND sky130_fd_pr__pfet_01v8_6KFL8S
C0 WL BL_IN 0.11791f
C1 GND BL_IN 0.11225f
C2 BL_NIN WL 0.06023f
C3 BL_N VDD 0.04917f
C4 BL_NIN GND 0.0643f
C5 VDD BL_IN 0.21734f
C6 BL_NIN VDD 0.1729f
C7 WL GND 0.04765f
C8 WL VDD 0.36318f
C9 VDD GND 0.15978f
C10 BL_N BL 0
C11 BL BL_IN 0.0109f
C12 BL_NIN BL 0.00177f
C13 BL WL 0.08926f
C14 BL GND 0.00163f
C15 BL VDD 0.81625f
C16 BL_N BL_IN 0.03664f
C17 BL_N BL_NIN 0.04099f
C18 BL_NIN BL_IN 0.07337f
C19 BL_N WL 0.09632f
C20 BL_N GND 0.06251f
C21 VDD 0 3.02205f
C22 BL_NIN 0 0.45842f
C23 GND 0 0.1696f
C24 BL_IN 0 0.41809f
C25 BL 0 0.63429f
C26 WL 0 1.19711f
C27 BL_N 0 1.11512f
.ends

