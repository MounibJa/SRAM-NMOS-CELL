magic
tech sky130A
magscale 1 2
timestamp 1764564536
<< error_s >>
rect 140 -300 380 -298
<< pwell >>
rect -180 320 620 440
rect -341 179 620 320
rect -180 100 620 179
<< psubdiff >>
rect -330 280 -220 310
rect -330 230 -300 280
rect -250 230 -220 280
rect -330 200 -220 230
<< psubdiffcont >>
rect -300 230 -250 280
<< locali >>
rect -320 280 -230 300
rect -320 230 -300 280
rect -250 230 -230 280
rect -320 210 -230 230
<< viali >>
rect 492 862 526 916
rect -300 230 -250 280
rect 492 -390 526 -350
<< metal1 >>
rect -440 400 -360 1040
rect 471 916 544 942
rect 130 820 160 880
rect 340 820 390 880
rect 471 862 492 916
rect 526 862 544 916
rect 630 870 710 1040
rect 471 853 544 862
rect 130 810 390 820
rect 374 772 420 776
rect 489 772 526 853
rect 629 820 710 870
rect 630 772 710 820
rect 0 700 120 760
rect 0 690 80 700
rect 374 697 711 772
rect 0 530 40 690
rect 374 688 420 697
rect 0 490 380 530
rect -90 440 0 450
rect -440 360 -140 400
rect -90 380 -80 440
rect -10 380 0 440
rect 340 380 380 490
rect -90 370 0 380
rect -440 -530 -360 360
rect -180 340 -140 360
rect 220 350 380 380
rect 450 430 540 440
rect 450 370 460 430
rect 530 370 540 430
rect -320 282 -230 300
rect -320 230 -302 282
rect -250 230 -230 282
rect -180 280 -80 340
rect 100 300 140 340
rect 340 300 380 350
rect 530 310 600 320
rect 0 250 140 300
rect -320 210 -230 230
rect 100 160 140 250
rect 184 290 290 300
rect 184 230 190 290
rect 280 230 290 290
rect 184 220 290 230
rect 340 250 460 300
rect 340 180 380 250
rect 530 220 540 310
rect 592 220 600 310
rect 530 200 600 220
rect 100 120 280 160
rect 100 50 160 120
rect 10 0 160 50
rect 10 -160 60 0
rect 10 -170 80 -160
rect 630 -169 710 697
rect 770 310 850 1040
rect 770 250 780 310
rect 840 250 850 310
rect 10 -240 120 -170
rect 379 -238 711 -169
rect 130 -300 390 -290
rect 130 -350 140 -300
rect 380 -350 390 -300
rect 481 -340 710 -238
rect 481 -348 540 -340
rect 130 -360 390 -350
rect 480 -350 540 -348
rect 480 -390 492 -350
rect 526 -390 540 -350
rect 480 -400 540 -390
rect 630 -529 710 -340
rect 770 -530 850 250
<< via1 >>
rect 160 820 340 880
rect -80 380 -10 440
rect 460 370 530 430
rect -302 280 -250 282
rect -302 230 -300 280
rect -300 230 -250 280
rect 190 230 280 290
rect 540 220 592 310
rect 780 250 840 310
rect 140 -350 380 -300
<< metal2 >>
rect -300 870 -230 1040
rect 130 870 160 880
rect -300 820 160 870
rect 340 820 390 880
rect -300 770 -230 820
rect 130 810 390 820
rect -300 690 -229 770
rect -300 290 -230 690
rect -90 440 0 450
rect -90 380 -80 440
rect -10 380 0 440
rect -90 370 0 380
rect 450 430 540 440
rect 450 370 460 430
rect 530 370 540 430
rect 450 360 540 370
rect 530 310 600 320
rect -320 282 -230 290
rect -320 230 -302 282
rect -250 270 -230 282
rect 180 290 290 300
rect 180 270 190 290
rect -250 240 190 270
rect -250 230 -230 240
rect -320 220 -230 230
rect 180 230 190 240
rect 280 230 290 290
rect 180 220 290 230
rect 530 220 540 310
rect 592 300 600 310
rect 770 310 850 320
rect 770 300 780 310
rect 592 250 780 300
rect 840 250 850 310
rect 592 240 850 250
rect 592 220 600 240
rect -300 -300 -230 220
rect 530 210 600 220
rect 130 -300 390 -290
rect -300 -350 140 -300
rect 380 -350 390 -300
rect -300 -530 -230 -350
rect 130 -360 390 -350
<< via2 >>
rect -80 380 -10 440
rect 460 370 530 430
<< metal3 >>
rect -560 440 920 450
rect -560 390 -80 440
rect -90 380 -80 390
rect -10 430 920 440
rect -10 390 460 430
rect -10 380 0 390
rect -90 370 0 380
rect 450 370 460 390
rect 530 390 920 430
rect 530 370 540 390
rect 450 360 540 370
use sky130_fd_pr__nfet_01v8_BHJCXL  sky130_fd_pr__nfet_01v8_BHJCXL_0
timestamp 1764448333
transform 0 1 238 -1 0 257
box -137 -138 137 138
use sky130_fd_pr__nfet_01v8_HKHAX8  sky130_fd_pr__nfet_01v8_HKHAX8_0
timestamp 1764459837
transform 1 0 -45 0 1 263
box -83 -163 83 163
use sky130_fd_pr__nfet_01v8_HKHAX8  sky130_fd_pr__nfet_01v8_HKHAX8_1
timestamp 1764459837
transform 1 0 491 0 1 261
box -83 -163 83 163
use sky130_fd_pr__pfet_01v8_6KFL8S  sky130_fd_pr__pfet_01v8_6KFL8S_0
timestamp 1764564536
transform -1 0 246 0 -1 731
box -316 -261 316 261
use sky130_fd_pr__pfet_01v8_6KFL8S  sky130_fd_pr__pfet_01v8_6KFL8S_1
timestamp 1764564536
transform 1 0 246 0 1 -209
box -316 -261 316 261
<< labels >>
rlabel metal1 654 1008 654 1008 1 VDD
port 1 n
rlabel metal1 778 1012 778 1012 1 BL
port 4 n
rlabel metal1 -412 994 -412 994 1 BL_N
port 5 n
rlabel metal2 -268 998 -268 998 1 GND
port 2 n
rlabel metal3 -520 418 -520 418 7 WL
port 3 w
rlabel metal1 360 316 360 316 1 BL_IN
port 6 n
rlabel metal1 126 150 126 150 5 BL_NIN
port 7 s
<< end >>
