magic
tech sky130A
magscale 1 2
timestamp 1764558790
<< pwell >>
rect 699 590 1479 930
rect 10 484 160 550
rect -194 110 660 484
<< psubdiff >>
rect 30 500 140 530
rect 30 450 60 500
rect 110 450 140 500
rect 30 420 140 450
<< psubdiffcont >>
rect 60 450 110 500
<< locali >>
rect 40 500 130 520
rect 40 450 60 500
rect 110 450 130 500
rect 40 430 130 450
<< viali >>
rect -900 654 -866 700
rect -900 620 -840 654
rect 60 450 110 500
rect -900 13 -820 50
rect -900 -20 -860 13
<< metal1 >>
rect -1100 300 -1000 1700
rect -700 1260 -380 1460
rect -20 1400 620 1480
rect -720 920 -400 1120
rect -180 1100 140 1300
rect 360 1100 680 1300
rect 920 1260 1240 1460
rect -920 700 -820 720
rect -920 620 -900 700
rect -920 600 -820 620
rect -720 680 -420 800
rect -180 760 140 960
rect 340 799 660 960
rect 900 940 1220 1140
rect 1500 820 1620 1700
rect 340 760 479 799
rect 645 760 660 799
rect 880 740 1620 820
rect -720 560 420 680
rect 40 502 130 520
rect 40 450 60 502
rect 112 450 130 502
rect 40 430 130 450
rect 340 380 420 560
rect 220 350 420 380
rect 340 346 420 350
rect 100 300 140 340
rect 340 300 418 346
rect -1100 240 -100 300
rect 0 250 140 300
rect -1100 -1040 -1000 240
rect -90 162 -10 180
rect -90 150 -80 162
rect -100 110 -80 150
rect -28 110 -10 162
rect 60 160 140 250
rect 184 290 290 300
rect 184 230 190 290
rect 280 230 290 290
rect 184 220 290 230
rect 340 250 480 300
rect 580 280 1120 300
rect 580 250 1040 280
rect 340 180 380 250
rect 590 240 1040 250
rect 1020 200 1040 240
rect 1100 200 1120 280
rect 1020 180 1120 200
rect -100 100 -10 110
rect 40 120 280 160
rect 490 152 570 160
rect -920 60 -800 80
rect -920 -20 -900 60
rect -820 -20 -800 60
rect -920 -40 -800 -20
rect -720 -300 -380 -100
rect 40 -140 160 120
rect 490 100 500 152
rect 560 100 570 152
rect 1500 -80 1620 740
rect -720 -620 -380 -420
rect -160 -460 180 -260
rect 340 -300 680 -100
rect 860 -140 1620 -80
rect -200 -740 140 -600
rect 340 -620 680 -420
rect 900 -460 1240 -260
rect -200 -800 660 -740
rect 880 -800 1220 -600
rect -160 -820 660 -800
rect 1500 -1040 1620 -140
rect 1700 260 1800 1700
rect 1700 200 1720 260
rect 1780 200 1800 260
rect 1700 -1040 1800 200
<< via1 >>
rect -900 654 -866 700
rect -866 654 -820 700
rect -900 620 -840 654
rect -840 620 -820 654
rect 60 500 112 502
rect 60 450 110 500
rect 110 450 112 500
rect -80 110 -28 162
rect 190 230 280 290
rect 1040 200 1100 280
rect -900 50 -820 60
rect -900 13 -820 50
rect -900 -20 -860 13
rect -860 -20 -820 13
rect 500 100 560 152
rect 1720 200 1780 260
<< metal2 >>
rect -1340 520 -1240 1700
rect -920 700 -820 720
rect -920 620 -900 700
rect -920 600 -820 620
rect -900 520 -840 600
rect -1340 502 120 520
rect -1340 450 60 502
rect 112 450 120 502
rect -1340 440 120 450
rect -1340 -1040 -1240 440
rect -900 80 -840 440
rect 50 430 120 440
rect 70 270 100 430
rect 180 290 290 300
rect 180 270 190 290
rect 70 240 190 270
rect 180 230 190 240
rect 280 230 290 290
rect 180 220 290 230
rect 1020 280 1120 300
rect 1020 200 1040 280
rect 1100 260 1800 280
rect 1100 200 1720 260
rect 1780 200 1800 260
rect 1020 180 1120 200
rect 1700 180 1800 200
rect -90 166 -10 180
rect -90 110 -80 166
rect -24 110 -10 166
rect -90 100 -10 110
rect 490 160 580 170
rect 490 100 500 160
rect 570 100 580 160
rect 490 90 580 100
rect -920 60 -800 80
rect -920 -20 -900 60
rect -820 -20 -800 60
rect -920 -40 -800 -20
<< via2 >>
rect -80 162 -24 166
rect -80 110 -28 162
rect -28 110 -24 162
rect 500 152 570 160
rect 500 100 560 152
rect 560 100 570 152
<< metal3 >>
rect -1560 166 1970 180
rect -1560 120 -80 166
rect -100 110 -80 120
rect -24 160 1970 166
rect -24 120 500 160
rect -24 110 -10 120
rect -100 90 -10 110
rect 480 100 500 120
rect 570 120 1970 160
rect 570 100 600 120
rect 480 80 600 100
use sky130_fd_pr__nfet_01v8_BHJCXL  sky130_fd_pr__nfet_01v8_BHJCXL_0
timestamp 1764448333
transform 0 1 238 -1 0 257
box -137 -138 137 138
use sky130_fd_pr__nfet_01v8_HKHAX8  sky130_fd_pr__nfet_01v8_HKHAX8_0
timestamp 1764459837
transform 1 0 533 0 1 283
box -83 -163 83 163
use sky130_fd_pr__nfet_01v8_HKHAX8  sky130_fd_pr__nfet_01v8_HKHAX8_1
timestamp 1764459837
transform 1 0 -57 0 1 283
box -83 -163 83 163
use sky130_fd_pr__res_xhigh_po_0p35_ZFXP64  sky130_fd_pr__res_xhigh_po_0p35_ZFXP64_0
timestamp 1764454615
transform 0 1 248 -1 0 1113
box -533 -1188 533 1188
use sky130_fd_pr__res_xhigh_po_0p35_ZFXP64  sky130_fd_pr__res_xhigh_po_0p35_ZFXP64_1
timestamp 1764454615
transform 0 -1 248 1 0 -447
box -533 -1188 533 1188
<< labels >>
rlabel metal1 1560 1660 1560 1660 1 VDD
port 1 n
rlabel metal1 1760 1660 1760 1660 1 BL
port 3 n
rlabel metal1 -1040 1660 -1040 1660 1 BL_N
port 4 n
rlabel metal2 -1300 1660 -1300 1660 1 GND
port 2 n
rlabel metal1 100 220 100 220 1 BL_NIN
port 6 n
rlabel metal1 380 300 380 300 1 BL_IN
port 5 n
rlabel metal3 -1500 150 -1500 150 7 WL
port 7 w
<< end >>
